`include "and64.v"
module and64_test;

reg signed [63:0] A, B;
wire signed [63:0] C;   
integer i;
output overflow;
reg [1:0] control;

and64 dut(.A(A), .B(B), .C(C),.overflow(overflow),.control(control));

initial begin
    
    $dumpfile("and64_test.vcd");
    $dumpvars(0,and64_test);

    A = 64'b0; B = 64'b0;

    $monitor("A = %b\nb = %b\nc = %b\n\n" , A, B, C);

    #100
    A = 64'b1111111111111111111111111111111111111111111111111111111111110000;
    B = 64'b1111111111111111111111111111111111111111111111111111111111111111;

    #100
    A = 64'b1111111111011111111111011111111111111111111111111111111111110000;
    B = 64'b1111111111011111111111011111111111111110111111111111111111111111;

    #100
    A = 64'b0111111111111111111111111111011111111111111111111111111111110000;
    B = 64'b1111111111111111111101111111111111111111111110111111111111111111;

end 
endmodule
